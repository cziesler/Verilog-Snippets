//===========================================================================//
// File name: tb_half_adder.v
// Author:    Cody Cziesler
//
// Description: Test bench for testing tb_half_adder.v
//
//===========================================================================//

module tb_half_adder ();

//---------------------------------------------------------------------------//
// Inputs to UUT
//---------------------------------------------------------------------------//
reg a;
reg b;

//---------------------------------------------------------------------------//
// Outputs from UUT
//---------------------------------------------------------------------------//
wire sum;
wire c_out;

//---------------------------------------------------------------------------//
// A lcv
//---------------------------------------------------------------------------//
integer i;

//---------------------------------------------------------------------------//
// Create the vpd file
//---------------------------------------------------------------------------//
initial begin
  $vcdpluson(tb_half_adder);
end

//---------------------------------------------------------------------------//
// Initialize signals and perform test
//---------------------------------------------------------------------------//
initial begin
  $display ("======================================");
  $display ("Starting tb_half_adder");

  for (i = 32'd0; i < 32'h4; i = i + 1) begin
    {a, b} = i;
    #1;
    if ( {c_out, sum} !== add (a, b) ) begin
      $display("ERROR - a[%b] + b[%b] !== c_out[%b], sum[%b] @ %0t",
        a, b, c_out, sum, $time);
    end
  end

  $display ("======================================");
  $finish ();
end

//---------------------------------------------------------------------------//
// UUT (half_adder.v)
//---------------------------------------------------------------------------//
half_adder half_adder_0 (
  .a(a),
  .b(b),
  .sum(sum),
  .c_out(c_out)
);

//---------------------------------------------------------------------------//
// Add two numbers
//---------------------------------------------------------------------------//
function [1:0] add;
  input a;
  input b;
begin
  add[1:0] = a + b;
end
endfunction

endmodule
